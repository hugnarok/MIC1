library verilog;
use verilog.vl_types.all;
entity MIC1_vlg_check_tst is
    port(
        O0              : in     vl_logic;
        O1              : in     vl_logic;
        O2              : in     vl_logic;
        O3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MIC1_vlg_check_tst;
